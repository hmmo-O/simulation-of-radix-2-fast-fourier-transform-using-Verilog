// Module Name: or31
module or31(a1,a2,a3,z );
input a1;
input a2;
input a3;
output z;
wire z;
assign z=a1|a2|a3;
endmodule