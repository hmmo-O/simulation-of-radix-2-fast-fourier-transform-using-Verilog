// Module Name: xor21
module xor21(a1,a2,z);
input a1;
input a2;
wire z;
output z;
assign z=a1^a2;
endmodule