// Module Name: or21
module or21(a1,a2,z );
input a1;
input a2;
output z;
assign z=a1|a2;
endmodule