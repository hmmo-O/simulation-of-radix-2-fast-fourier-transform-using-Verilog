// Module name: and21
module and21(a1,a2,z );
input a1;
input a2;
output z;
wire z;
assign z=a1&a2;
endmodule