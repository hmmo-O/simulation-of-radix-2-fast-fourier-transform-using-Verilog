// Module name: and31
module and31(a1,a2,a3,z );
input a1;
input a2;
input a3;
output z;

wire z;
assign z=a1&a2&a3;
endmodule