// Module Name: and41
module and41(a1,a2,a3,z,a4 );
input a1;
input a2;
input a3;
input a4;
output z;
wire z;
assign z=a1&a2&a3&a4;
endmodule